/* $Author: sinclair $ */
/* $LastChangedDate: 2020-02-09 17:03:45 -0600 (Sun, 09 Feb 2020) $ */
/* $Rev: 46 $ */
module proc (/*AUTOARG*/
    // Outputs
        err, 
    // Inputs
    clk, rst
    );

    input clk;
    input rst;

    output err;

    // None of the above lines can be modified

    // OR all the err ouputs for every sub-module and assign it as this
    // err output
    
    // As desribed in the homeworks, use the err signal to trap corner
    // cases that you think are illegal in your statemachines
    
    
    /* your code here -- should include instantiations of fetch, decode, execute, mem and wb modules */
    
    wire RegDst, Jump, Branch, MemRead, MemToReg, MemWrite, ALU_Src, RegWrite; 
    wire [4:0] ALU_op;
    wire control_err;
    wire halt;
    wire five_bit_imm;
    wire ZeroExtend;
    wire alu_ofl;

    //write_back Outputs
    wire [15:0] wb_out; 
    wire [15:0] wb_pc;

    //data_mem Outputs
    wire [15:0] branch_or_pc;
    wire [15:0] data_mem_out;

    //ALU Outputs
    wire [15:0] ALU_result;
    wire zero;
    wire [15:0] branch_result;
    wire alu_err;
    wire ltz;
    wire [15:0] jump_out;

    //Decode Outputs
    wire [15:0] jumpAddr;
    wire [15:0] read1data;
    wire [15:0] read2data;
    wire [15:0] immediate;
    wire decode_err;

    //Fetch Outputs
    wire [15:0] next_pc;
    wire [15:0] instruction;
    wire fetch_err;

    //ALU Control Outputs
    wire [2:0] op_to_alu;
    wire invA, invB;
    wire sign;
    wire cin;
    wire passA;
    wire passB;

    
    fetch fetch0(//Input
                        .pc(wb_pc), .clk(clk), .rst(rst), 
                        //Outputs
                        .next_pc(next_pc), .instr(instruction), .err(fetch_err));

    decode decode0(//Inputs
                        .instruction(instruction), .RegWrite(RegWrite), .RegDst(RegDst), .writeData(wb_out),
                        .clk(clk), .rst(rst), .pc(next_pc[15:0]), .five_bit_imm(five_bit_imm), .ZeroExtend(ZeroExtend),
                        .MemWrite(MemWrite),
                        //Outputs
                        .jumpAddr(jumpAddr), .read1data(read1data), .read2data(read2data), .immediate(immediate),
                        .err(decode_err));  
    
    
    execute exec0 ( //Inputs
                        .alu_op(op_to_alu), .ALUSrc(ALU_Src), .read1data(read1data), .read2data(read2data), 
                        .immediate(immediate), .pc(next_pc), .invA(invA), .invB(invB), .cin(cin), .sign(sign),  
                        .passThroughA(passA), .passThroughB(passB), .instr_op(ALU_op), .MemWrite(MemWrite),
                        .jump_in(jumpAddr),
                        //Outputs
                        .ALU_result(ALU_result), .branch_result(branch_result), .zero(zero), .err(alu_err),
                        .ltz(ltz), .jump_out(jump_out));  
    
    
    data_mem memory0(.memWrite(MemWrite), .memRead(MemRead), .ALU_result(ALU_result), .writedata(read2data), 
                    .readData(data_mem_out), .zero(zero), .Branch(Branch), .branchAddr(branch_result), .pc(next_pc), 
                    .halt(halt), .ltz(ltz), .branch_op(ALU_op[1:0]), .branch_or_pc(branch_or_pc), .clk(clk), .rst(rst));  
    
    
    wb wb0 (.mem_data(data_mem_out), .ALU_result(ALU_result), .MemToReg(MemToReg), .jumpAddr(jump_out), 
                    .branch_or_pc(branch_or_pc), .Jump(Jump), .pc(wb_pc), .out_data(wb_out)); 
    
    
    control control0( //Inputs
                        .instruction_op(instruction[15:11]),
                        //Outputs 
                        .RegDst(RegDst), .Jump(Jump), .Branch(Branch), .MemRead(MemRead), .MemToReg(MemToReg), .halt(halt),
                        .ALU_op(ALU_op), .MemWrite(MemWrite), .ALUSrc(ALU_Src), .RegWrite(RegWrite), .err(control_err),
                        .five_bit_imm(five_bit_imm), .ZeroExtend(ZeroExtend));

    alu_control actl0(//Inputs
                        .ALU_op(ALU_op), .ALU_funct(instruction[1:0]), 
                        //Outputs
                        .invA(invA), .invB(invB), .op_to_alu(op_to_alu), .cin(cin), .sign(sign), .passA(passA), .passB(passB));
endmodule // proc
// DUMMY LINE FOR REV CONTROL :0:
