module forward_mem(/* input */ 
    /* output */  );
    
endmodule
