module forward_mem(/* input */ MemWriteExMem, 
    /* output */  );
    
endmodule
